////////////////////////////////////////////////////////////////////////////////
//
// Filename: 	rtcbare.v
//
// Project:	A Wishbone Controlled Real--time Clock Core, w/ GPS synch
//
// Purpose:	This is the bare RTC clock logic.
//
// Creator:	Dan Gisselquist, Ph.D.
//		Gisselquist Technology, LLC
//
////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2015-2018, Gisselquist Technology, LLC
//
// This program is free software (firmware): you can redistribute it and/or
// modify it under the terms of  the GNU General Public License as published
// by the Free Software Foundation, either version 3 of the License, or (at
// your option) any later version.
//
// This program is distributed in the hope that it will be useful, but WITHOUT
// ANY WARRANTY; without even the implied warranty of MERCHANTIBILITY or
// FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
// for more details.
//
// You should have received a copy of the GNU General Public License along
// with this program.  (It's in the $(ROOT)/doc directory.  Run make with no
// target there if the PDF file isn't present.)  If not, see
// <http://www.gnu.org/licenses/> for a copy.
//
// License:	GPL, v3, as defined and found on www.gnu.org,
//		http://www.gnu.org/licenses/gpl.html
//
//
////////////////////////////////////////////////////////////////////////////////
//
//
`default_nettype	none
//
module	rtcbare(i_clk, i_reset,
		// Wishbone interface
		i_pps, i_wr, i_data, i_valid,
		// Output registers
		o_data, // multiplexed based upon i_wb_addr
		// A once-per-day strobe on the last clock of the day
		o_ppd);
	//
	input	wire		i_clk, i_reset;
	//
	input	wire		i_pps, i_wr;
	input	wire	[21:0]	i_data;
	input	wire	[2:0]	i_valid;
	output	wire	[21:0]	o_data;
	output	wire		o_ppd;

	reg	[21:0]	bcd_clock, next_clock;
	reg	[5:0]	carry;
	reg		pre_ppd;

	initial	pre_ppd = 1'b0;
	always @(posedge i_clk)
	if (i_reset)
		pre_ppd <= 1'b0;
	else
		pre_ppd <= (bcd_clock == 22'h23_59_59);

	initial	next_clock = 22'h00_00_01;
	always @(posedge i_clk)
	if (i_reset)
		next_clock <= 22'h00_00_01;
	else begin
		// Takes 7 clocks to converge

		// Seconds
		carry[0] <= (bcd_clock[ 3: 0] >=  4'h9);
		carry[1] <= (bcd_clock[ 7: 4] >=  4'h5)&&( carry[  0]);
		// Minutes
		carry[2] <= (bcd_clock[11: 8] >=  4'h9)&&(&carry[1:0]);
		carry[3] <= (bcd_clock[15:12] >=  4'h5)&&(&carry[2:0]);
		// Hours
		carry[4] <= (bcd_clock[19:16] >=  4'h9)&&(&carry[3:0]);
		carry[5] <= (bcd_clock[21:16] >= 6'h23)&&(&carry[3:0]);

		// Seconds
		if (carry[0])
			next_clock[3:0] <= 4'h0;
		else
			next_clock[3:0] <= bcd_clock[3:0] + 4'h1;

		if (carry[1])
			next_clock[7:4] <= 4'h0;
		else if (carry[0])
			next_clock[7:4] <= bcd_clock[7:4] + 4'h1;
		else
			next_clock[7:4] <= bcd_clock[7:4];

		// Minutes
		if (carry[2])
			next_clock[11:8] <= 4'h0;
		else if (carry[1])
			next_clock[11:8] <= bcd_clock[11:8] + 4'h1;
		else
			next_clock[11:8] <= bcd_clock[11:8];

		if (carry[3])
			next_clock[15:12] <= 4'h0;
		else if (carry[2])
			next_clock[15:12] <= bcd_clock[15:12] + 4'h1;
		else
			next_clock[15:12] <= bcd_clock[15:12];

		// Hours
		if ((carry[4])||(carry[5]))
			next_clock[19:16] <= 4'h0;
		else if (carry[3])
			next_clock[19:16] <= bcd_clock[19:16] + 4'h1;
		else
			next_clock[19:16] <= bcd_clock[19:16];

		if (carry[5])
			next_clock[21:20] <= 2'h0;
		else if (carry[4])
			next_clock[21:20] <= bcd_clock[21:20] + 2'h1;
		else
			next_clock[21:20] <= bcd_clock[21:20];
	end

	reg	[2:0]	suppressed, suppress_count;

	initial	suppressed = 3'h7;
	initial	suppress_count = 3'h5;
	always @(posedge i_clk)
	if (i_reset)
	begin
		suppressed <= 3'h7;
		suppress_count <= 3'h5;
	end else if ((i_wr)&&(|i_valid))
	begin
		suppressed[0] <= (suppressed[0])||(i_valid[  0]!=1'b0);
		suppressed[1] <= (suppressed[1])||(i_valid[1:0]!=2'b00);
		suppressed[2] <= (suppressed[2])||(i_valid[2:0]!=3'b000);
		suppress_count <= 3'h5;
	end else if (suppress_count > 0)
		suppress_count <= suppress_count - 1;
	else
		suppressed <= 0;

	initial	bcd_clock = 0;
	always @(posedge i_clk)
	if (i_reset)
		bcd_clock <= 0;
	else begin
		if (i_pps)
		begin
			if (!suppressed[0])
				bcd_clock[7:0] <= next_clock[7:0];
			if (!suppressed[1])
				bcd_clock[15:8] <= next_clock[15:8];
			if (!suppressed[2])
				bcd_clock[21:16] <= next_clock[21:16];
		end
		if ((i_wr)&&(i_valid[0]))
			bcd_clock[7:0] <= i_data[7:0];
		if ((i_wr)&&(i_valid[1]))
			bcd_clock[15:8] <= i_data[15:8];
		if ((i_wr)&&(i_valid[2]))
			bcd_clock[21:16] <= i_data[21:16];
	end

	assign	o_data = bcd_clock;
	assign	o_ppd  = (pre_ppd)&&(i_pps);

`ifdef	FORMAL
`ifdef	RTCBARE
`define	ASSUME	assume
`define	ASSERT	assert
`else
`define	ASSUME	assert
`define	ASSERT	assume
`endif

	reg	f_past_valid;
	initial	f_past_valid = 1'b0;
	always @(posedge i_clk)
		f_past_valid <= 1'b1;

	//
	always @(*)
	begin
		`ASSERT(bcd_clock[ 3: 0] <= 4'h9);
		`ASSERT(bcd_clock[ 7: 4] <= 4'h5);
		`ASSERT(bcd_clock[11: 8] <= 4'h9);
		`ASSERT(bcd_clock[15:12] <= 4'h5);
		`ASSERT(bcd_clock[19:16] <= 4'h9);
		`ASSERT(bcd_clock[21:16] <= 6'h23);
	end


	always @(*)
	if (i_wr)
	begin
		if (i_valid[0])
		begin
			`ASSUME(i_data[ 3: 0] <= 4'h9);
			`ASSUME(i_data[ 7: 4] <= 4'h5);
		end

		if (i_valid[1])
		begin
			`ASSUME(i_data[11: 8] <= 4'h9);
			`ASSUME(i_data[15:12] <= 4'h5);
		end

		if (i_valid[2])
		begin
			`ASSUME(i_data[19:16] <= 4'h9);
			`ASSUME(i_data[21:16] <= 8'h23);
		end
	end

	always @(*)
	begin
		`ASSERT(bcd_clock[ 3: 0] <= 4'h9);
		`ASSERT(bcd_clock[ 7: 4] <= 4'h5);
		`ASSERT(bcd_clock[11: 8] <= 4'h9);
		`ASSERT(bcd_clock[15:12] <= 4'h5);
		`ASSERT(bcd_clock[19:16] <= 4'h9);
		`ASSERT(bcd_clock[21:16] <= 8'h23);
	end

	reg	[7:0]	f_past_pps;
	initial	f_past_pps = 0;
	always @(posedge i_clk)
	if (i_reset)
		f_past_pps <= 0;
	else if (i_pps)
		f_past_pps <= 8'hff;
	else
		f_past_pps <= { f_past_pps[6:0], 1'b0 };

	always @(*)
	if (f_past_pps[7])
		`ASSUME(!i_pps);

	always @(*)
		`ASSERT(suppress_count <= 3'h5);
	always @(*)
	if (suppressed[0])
		`ASSERT(suppressed[1]);
	always @(*)
	if (suppressed[1])
		`ASSERT(suppressed[2]);


`endif
endmodule
